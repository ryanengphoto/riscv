`timescale 1ns / 1ps
// =============================================================================
// ChaCha20 Full Block Testbench
// =============================================================================
// Dedicated testbench for running the complete ChaCha20 block algorithm.
// Features:
//   - Large instruction memory (256 words)
//   - Large data memory (1024 words)
//   - ChaCha20 RFC 7539 test vectors
// =============================================================================

`include "common_tasks.svh"

module tb_chacha20();

    // =========================================================================
    // Test Statistics
    // =========================================================================
    static int checked, errors;

    // =========================================================================
    // DUT Interface Signals
    // =========================================================================
    logic clk;
    logic rst;
    logic [31:0] imem_addr;
    logic [31:0] imem_data;
    logic dmem_read;
    logic dmem_write;
    logic [31:0] dmem_addr;
    logic [31:0] dmem_wdata;
    logic [31:0] dmem_rdata;

    // =========================================================================
    // Memory Models (LARGER for ChaCha20)
    // =========================================================================
    
    // Instruction memory (256 words = 1KB)
    logic [31:0] instruction_mem [0:255];
    
    // Data memory (1024 words = 4KB)
    logic [31:0] data_mem [0:1023];
    
    // Initialize memories
    initial begin
        for (int i = 0; i < 256; i++) begin
            instruction_mem[i] = 32'h00000013; // ADDI x0, x0, 0 (NOP)
        end
        for (int i = 0; i < 1024; i++) begin
            data_mem[i] = 32'h0;
        end
    end

    // Instruction memory read (combinational)
    always_comb begin
        if (imem_addr[31:2] < 256) begin
            imem_data = instruction_mem[imem_addr[31:2]];
        end else begin
            imem_data = 32'h00000013; // NOP for out-of-range
        end
    end

    // Data memory write (synchronous)
    always_ff @(posedge clk) begin
        if (dmem_write && (dmem_addr[31:2] < 1024)) begin
            data_mem[dmem_addr[31:2]] <= dmem_wdata;
        end
    end

    // Data memory read (combinational)
    always_comb begin
        if (dmem_read && (dmem_addr[31:2] < 1024)) begin
            dmem_rdata = data_mem[dmem_addr[31:2]];
        end else begin
            dmem_rdata = 32'h0;
        end
    end

    // =========================================================================
    // DUT Instantiation
    // =========================================================================
    riscv_cpu u_riscv_cpu (
        .clk(clk),
        .rst(rst),
        .imem_addr(imem_addr),
        .imem_data(imem_data),
        .dmem_read(dmem_read),
        .dmem_write(dmem_write),
        .dmem_addr(dmem_addr),
        .dmem_wdata(dmem_wdata),
        .dmem_rdata(dmem_rdata)
    );

    // =========================================================================
    // Clock Generation
    // =========================================================================
    initial clk = 1'b0;
    always #5 clk = ~clk;  // 100MHz clock (10ns period)

    // =========================================================================
    // ChaCha20 Test Vector (RFC 7539)
    // =========================================================================
    task automatic load_chacha20_test_vector();
        // ChaCha20 Input State:
        // Constants: "expand 32-byte k"
        data_mem[0]  = 32'h61707865;  // "expa"
        data_mem[1]  = 32'h3320646e;  // "nd 3"
        data_mem[2]  = 32'h79622d32;  // "2-by"
        data_mem[3]  = 32'h6b206574;  // "te k"
        
        // Key (256 bits = 8 words) - Non-zero key for testing
        data_mem[4]  = 32'h03020100;  // Key word 0
        data_mem[5]  = 32'h07060504;  // Key word 1
        data_mem[6]  = 32'h0b0a0908;  // Key word 2
        data_mem[7]  = 32'h0f0e0d0c;  // Key word 3
        data_mem[8]  = 32'h13121110;  // Key word 4
        data_mem[9]  = 32'h17161514;  // Key word 5
        data_mem[10] = 32'h1b1a1918;  // Key word 6
        data_mem[11] = 32'h1f1e1d1c;  // Key word 7
        
        // Counter (32 bits)
        data_mem[12] = 32'h00000001;
        
        // Nonce (96 bits = 3 words) - Non-zero nonce
        data_mem[13] = 32'h09000000;  // Nonce word 0
        data_mem[14] = 32'h4a000000;  // Nonce word 1
        data_mem[15] = 32'h00000000;  // Nonce word 2
    endtask

    // =========================================================================
    // Load Assembled ChaCha20 Program
    // Generated by: python3 tools/rv32_assembler.py sim/asm/chacha20_full.s
    // =========================================================================
    task automatic load_chacha20_program();
        instruction_mem[0] = 32'h00000137;  // lui     sp, 0
        instruction_mem[1] = 32'h1FC10113;  // addi    sp, sp, 0x1FC
        instruction_mem[2] = 32'h00000F13;  // addi    t5, x0, 0
        instruction_mem[3] = 32'h04000513;  // addi    a0, x0, 0x40
        instruction_mem[4] = 32'h00000593;  // addi    a1, x0, 0x00
        instruction_mem[5] = 32'h00C0006F;  // j       12
        instruction_mem[6] = 32'h00100F93;  // addi    t6, x0, 1
        instruction_mem[7] = 32'h21F02223;  // sw      t6, 0x204(x0)
        instruction_mem[8] = 32'h00000013;  // nop
        instruction_mem[9] = 32'h00000293;  // addi    t0, x0, 0
        instruction_mem[10] = 32'h01000313;  // addi    t1, x0, 16
        instruction_mem[11] = 32'h08000393;  // addi    t2, x0, 0x80
        instruction_mem[12] = 32'h0005AE03;  // lw      t3, 0(a1)
        instruction_mem[13] = 32'h01C3A023;  // sw      t3, 0(t2)
        instruction_mem[14] = 32'h00458593;  // addi    a1, a1, 4
        instruction_mem[15] = 32'h00438393;  // addi    t2, t2, 4
        instruction_mem[16] = 32'h00128293;  // addi    t0, t0, 1
        instruction_mem[17] = 32'hFE62C6E3;  // blt     t0, t1, -20
        instruction_mem[18] = 32'h00000593;  // addi    a1, x0, 0x00
        instruction_mem[19] = 32'h08000393;  // addi    t2, x0, 0x80
        instruction_mem[20] = 32'h0003A403;  // lw      s0, 0(t2)
        instruction_mem[21] = 32'h0043A483;  // lw      s1, 4(t2)
        instruction_mem[22] = 32'h0083A903;  // lw      s2, 8(t2)
        instruction_mem[23] = 32'h00C3A983;  // lw      s3, 12(t2)
        instruction_mem[24] = 32'h0103AA03;  // lw      s4, 16(t2)
        instruction_mem[25] = 32'h0143AA83;  // lw      s5, 20(t2)
        instruction_mem[26] = 32'h0183AB03;  // lw      s6, 24(t2)
        instruction_mem[27] = 32'h01C3AB83;  // lw      s7, 28(t2)
        instruction_mem[28] = 32'h0203A603;  // lw      a2, 32(t2)
        instruction_mem[29] = 32'h0243A683;  // lw      a3, 36(t2)
        instruction_mem[30] = 32'h0283A703;  // lw      a4, 40(t2)
        instruction_mem[31] = 32'h02C3A783;  // lw      a5, 44(t2)
        instruction_mem[32] = 32'h0303A803;  // lw      a6, 48(t2)
        instruction_mem[33] = 32'h0343A883;  // lw      a7, 52(t2)
        instruction_mem[34] = 32'h0383AE03;  // lw      t3, 56(t2)
        instruction_mem[35] = 32'h03C3AE83;  // lw      t4, 60(t2)
        instruction_mem[36] = 32'h00000293;  // addi    t0, x0, 0
        instruction_mem[37] = 32'h00A00313;  // addi    t1, x0, 10
        // === Column rounds ===
        instruction_mem[38] = 32'h01440433;  // add     s0, s0, s4
        instruction_mem[39] = 32'h00884833;  // xor     a6, a6, s0
        instruction_mem[40] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[41] = 32'h61F81833;  // rol     a6, a6, t6
        instruction_mem[42] = 32'h01060633;  // add     a2, a2, a6
        instruction_mem[43] = 32'h00C64A33;  // xor     s4, s4, a2
        instruction_mem[44] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[45] = 32'h61FA1A33;  // rol     s4, s4, t6
        instruction_mem[46] = 32'h01440433;  // add     s0, s0, s4
        instruction_mem[47] = 32'h00884833;  // xor     a6, a6, s0
        instruction_mem[48] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[49] = 32'h61F81833;  // rol     a6, a6, t6
        instruction_mem[50] = 32'h01060633;  // add     a2, a2, a6
        instruction_mem[51] = 32'h00C64A33;  // xor     s4, s4, a2
        instruction_mem[52] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[53] = 32'h61FA1A33;  // rol     s4, s4, t6
        instruction_mem[54] = 32'h015484B3;  // add     s1, s1, s5
        instruction_mem[55] = 32'h0098C8B3;  // xor     a7, a7, s1
        instruction_mem[56] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[57] = 32'h61F898B3;  // rol     a7, a7, t6
        instruction_mem[58] = 32'h011686B3;  // add     a3, a3, a7
        instruction_mem[59] = 32'h00D6CAB3;  // xor     s5, s5, a3
        instruction_mem[60] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[61] = 32'h61FA9AB3;  // rol     s5, s5, t6
        instruction_mem[62] = 32'h015484B3;  // add     s1, s1, s5
        instruction_mem[63] = 32'h0098C8B3;  // xor     a7, a7, s1
        instruction_mem[64] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[65] = 32'h61F898B3;  // rol     a7, a7, t6
        instruction_mem[66] = 32'h011686B3;  // add     a3, a3, a7
        instruction_mem[67] = 32'h00D6CAB3;  // xor     s5, s5, a3
        instruction_mem[68] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[69] = 32'h61FA9AB3;  // rol     s5, s5, t6
        instruction_mem[70] = 32'h01690933;  // add     s2, s2, s6
        instruction_mem[71] = 32'h012E4E33;  // xor     t3, t3, s2
        instruction_mem[72] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[73] = 32'h61FE1E33;  // rol     t3, t3, t6
        instruction_mem[74] = 32'h01C70733;  // add     a4, a4, t3
        instruction_mem[75] = 32'h00E74B33;  // xor     s6, s6, a4
        instruction_mem[76] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[77] = 32'h61FB1B33;  // rol     s6, s6, t6
        instruction_mem[78] = 32'h01690933;  // add     s2, s2, s6
        instruction_mem[79] = 32'h012E4E33;  // xor     t3, t3, s2
        instruction_mem[80] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[81] = 32'h61FE1E33;  // rol     t3, t3, t6
        instruction_mem[82] = 32'h01C70733;  // add     a4, a4, t3
        instruction_mem[83] = 32'h00E74B33;  // xor     s6, s6, a4
        instruction_mem[84] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[85] = 32'h61FB1B33;  // rol     s6, s6, t6
        instruction_mem[86] = 32'h017989B3;  // add     s3, s3, s7
        instruction_mem[87] = 32'h013ECEB3;  // xor     t4, t4, s3
        instruction_mem[88] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[89] = 32'h61FE9E33;  // rol     t4, t4, t6
        instruction_mem[90] = 32'h01D787B3;  // add     a5, a5, t4
        instruction_mem[91] = 32'h00F7CB33;  // xor     s7, s7, a5
        instruction_mem[92] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[93] = 32'h61FB9B33;  // rol     s7, s7, t6
        instruction_mem[94] = 32'h017989B3;  // add     s3, s3, s7
        instruction_mem[95] = 32'h013ECEB3;  // xor     t4, t4, s3
        instruction_mem[96] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[97] = 32'h61FE9E33;  // rol     t4, t4, t6
        instruction_mem[98] = 32'h01D787B3;  // add     a5, a5, t4
        instruction_mem[99] = 32'h00F7CB33;  // xor     s7, s7, a5
        instruction_mem[100] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[101] = 32'h61FB9B33;  // rol     s7, s7, t6
        // === Diagonal rounds ===
        instruction_mem[102] = 32'h01540433;  // add     s0, s0, s5
        instruction_mem[103] = 32'h008ECEB3;  // xor     t4, t4, s0
        instruction_mem[104] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[105] = 32'h61FE9E33;  // rol     t4, t4, t6
        instruction_mem[106] = 32'h01D70733;  // add     a4, a4, t4
        instruction_mem[107] = 32'h00E6CAB3;  // xor     s5, s5, a4
        instruction_mem[108] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[109] = 32'h61FA9AB3;  // rol     s5, s5, t6
        instruction_mem[110] = 32'h01540433;  // add     s0, s0, s5
        instruction_mem[111] = 32'h008ECEB3;  // xor     t4, t4, s0
        instruction_mem[112] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[113] = 32'h61FE9E33;  // rol     t4, t4, t6
        instruction_mem[114] = 32'h01D70733;  // add     a4, a4, t4
        instruction_mem[115] = 32'h00E6CAB3;  // xor     s5, s5, a4
        instruction_mem[116] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[117] = 32'h61FA9AB3;  // rol     s5, s5, t6
        instruction_mem[118] = 32'h016484B3;  // add     s1, s1, s6
        instruction_mem[119] = 32'h00984833;  // xor     a6, a6, s1
        instruction_mem[120] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[121] = 32'h61F81833;  // rol     a6, a6, t6
        instruction_mem[122] = 32'h010787B3;  // add     a5, a5, a6
        instruction_mem[123] = 32'h00F74B33;  // xor     s6, s6, a5
        instruction_mem[124] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[125] = 32'h61FB1B33;  // rol     s6, s6, t6
        instruction_mem[126] = 32'h016484B3;  // add     s1, s1, s6
        instruction_mem[127] = 32'h00984833;  // xor     a6, a6, s1
        instruction_mem[128] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[129] = 32'h61F81833;  // rol     a6, a6, t6
        instruction_mem[130] = 32'h010787B3;  // add     a5, a5, a6
        instruction_mem[131] = 32'h00F74B33;  // xor     s6, s6, a5
        instruction_mem[132] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[133] = 32'h61FB1B33;  // rol     s6, s6, t6
        instruction_mem[134] = 32'h01790933;  // add     s2, s2, s7
        instruction_mem[135] = 32'h0128C8B3;  // xor     a7, a7, s2
        instruction_mem[136] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[137] = 32'h61F898B3;  // rol     a7, a7, t6
        instruction_mem[138] = 32'h01160633;  // add     a2, a2, a7
        instruction_mem[139] = 32'h00C64B33;  // xor     s7, s7, a2
        instruction_mem[140] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[141] = 32'h61FB9B33;  // rol     s7, s7, t6
        instruction_mem[142] = 32'h01790933;  // add     s2, s2, s7
        instruction_mem[143] = 32'h0128C8B3;  // xor     a7, a7, s2
        instruction_mem[144] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[145] = 32'h61F898B3;  // rol     a7, a7, t6
        instruction_mem[146] = 32'h01160633;  // add     a2, a2, a7
        instruction_mem[147] = 32'h00C64B33;  // xor     s7, s7, a2
        instruction_mem[148] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[149] = 32'h61FB9B33;  // rol     s7, s7, t6
        instruction_mem[150] = 32'h014989B3;  // add     s3, s3, s4
        instruction_mem[151] = 32'h013E4E33;  // xor     t3, t3, s3
        instruction_mem[152] = 32'h01000F93;  // addi    t6, x0, 16
        instruction_mem[153] = 32'h61FE1E33;  // rol     t3, t3, t6
        instruction_mem[154] = 32'h01C686B3;  // add     a3, a3, t3
        instruction_mem[155] = 32'h00D64A33;  // xor     s4, s4, a3
        instruction_mem[156] = 32'h00C00F93;  // addi    t6, x0, 12
        instruction_mem[157] = 32'h61FA1A33;  // rol     s4, s4, t6
        instruction_mem[158] = 32'h014989B3;  // add     s3, s3, s4
        instruction_mem[159] = 32'h013E4E33;  // xor     t3, t3, s3
        instruction_mem[160] = 32'h00800F93;  // addi    t6, x0, 8
        instruction_mem[161] = 32'h61FE1E33;  // rol     t3, t3, t6
        instruction_mem[162] = 32'h01C686B3;  // add     a3, a3, t3
        instruction_mem[163] = 32'h00D64A33;  // xor     s4, s4, a3
        instruction_mem[164] = 32'h00700F93;  // addi    t6, x0, 7
        instruction_mem[165] = 32'h61FA1A33;  // rol     s4, s4, t6
        // Loop control
        instruction_mem[166] = 32'h00128293;  // addi    t0, t0, 1
        instruction_mem[167] = 32'hDE62CEE3;  // blt     t0, t1, -516
        // Add original state back
        instruction_mem[168] = 32'h00000393;  // addi    t2, x0, 0x00
        instruction_mem[169] = 32'h0003AF03;  // lw      t5, 0(t2)
        instruction_mem[170] = 32'h01E40433;  // add     s0, s0, t5
        instruction_mem[171] = 32'h0043AF03;  // lw      t5, 4(t2)
        instruction_mem[172] = 32'h01E484B3;  // add     s1, s1, t5
        instruction_mem[173] = 32'h0083AF03;  // lw      t5, 8(t2)
        instruction_mem[174] = 32'h01E90933;  // add     s2, s2, t5
        instruction_mem[175] = 32'h00C3AF03;  // lw      t5, 12(t2)
        instruction_mem[176] = 32'h01E989B3;  // add     s3, s3, t5
        instruction_mem[177] = 32'h0103AF03;  // lw      t5, 16(t2)
        instruction_mem[178] = 32'h01EA0A33;  // add     s4, s4, t5
        instruction_mem[179] = 32'h0143AF03;  // lw      t5, 20(t2)
        instruction_mem[180] = 32'h01EA8AB3;  // add     s5, s5, t5
        instruction_mem[181] = 32'h0183AF03;  // lw      t5, 24(t2)
        instruction_mem[182] = 32'h01EB0B33;  // add     s6, s6, t5
        instruction_mem[183] = 32'h01C3AF03;  // lw      t5, 28(t2)
        instruction_mem[184] = 32'h01EB8BB3;  // add     s7, s7, t5
        instruction_mem[185] = 32'h0203AF03;  // lw      t5, 32(t2)
        instruction_mem[186] = 32'h01E60633;  // add     a2, a2, t5
        instruction_mem[187] = 32'h0243AF03;  // lw      t5, 36(t2)
        instruction_mem[188] = 32'h01E686B3;  // add     a3, a3, t5
        instruction_mem[189] = 32'h0283AF03;  // lw      t5, 40(t2)
        instruction_mem[190] = 32'h01E70733;  // add     a4, a4, t5
        instruction_mem[191] = 32'h02C3AF03;  // lw      t5, 44(t2)
        instruction_mem[192] = 32'h01E787B3;  // add     a5, a5, t5
        instruction_mem[193] = 32'h0303AF03;  // lw      t5, 48(t2)
        instruction_mem[194] = 32'h01E80833;  // add     a6, a6, t5
        instruction_mem[195] = 32'h0343AF03;  // lw      t5, 52(t2)
        instruction_mem[196] = 32'h01E888B3;  // add     a7, a7, t5
        instruction_mem[197] = 32'h0383AF03;  // lw      t5, 56(t2)
        instruction_mem[198] = 32'h01EE0E33;  // add     t3, t3, t5
        instruction_mem[199] = 32'h03C3AF03;  // lw      t5, 60(t2)
        instruction_mem[200] = 32'h01EE8EB3;  // add     t4, t4, t5
        // Store output
        instruction_mem[201] = 32'h04802023;  // sw      s0, 0x40(x0)
        instruction_mem[202] = 32'h04902223;  // sw      s1, 0x44(x0)
        instruction_mem[203] = 32'h05202423;  // sw      s2, 0x48(x0)
        instruction_mem[204] = 32'h05302623;  // sw      s3, 0x4C(x0)
        instruction_mem[205] = 32'h05402823;  // sw      s4, 0x50(x0)
        instruction_mem[206] = 32'h05502A23;  // sw      s5, 0x54(x0)
        instruction_mem[207] = 32'h05602C23;  // sw      s6, 0x58(x0)
        instruction_mem[208] = 32'h05702E23;  // sw      s7, 0x5C(x0)
        instruction_mem[209] = 32'h06C02023;  // sw      a2, 0x60(x0)
        instruction_mem[210] = 32'h06D02223;  // sw      a3, 0x64(x0)
        instruction_mem[211] = 32'h06E02423;  // sw      a4, 0x68(x0)
        instruction_mem[212] = 32'h06F02623;  // sw      a5, 0x6C(x0)
        instruction_mem[213] = 32'h07002823;  // sw      a6, 0x70(x0)
        instruction_mem[214] = 32'h07102A23;  // sw      a7, 0x74(x0)
        instruction_mem[215] = 32'h07C02C23;  // sw      t3, 0x78(x0)
        instruction_mem[216] = 32'h07D02E23;  // sw      t4, 0x7C(x0)
        // Store round counter and integrity check
        instruction_mem[217] = 32'h20502023;  // sw      t0, 0x200(x0)
        instruction_mem[218] = 32'h60241F13;  // cpop    t5, s0 (I-type, correct RISC-V Zbb spec)
        instruction_mem[219] = 32'h21E02223;  // sw      t5, 0x204(x0)
        // Halt (infinite loop)
        instruction_mem[220] = 32'h00000013;  // nop
        instruction_mem[221] = 32'hFFDFF06F;  // j       -4 (halt loop)
    endtask

    // =========================================================================
    // Simple Loop Test (verify branch works)
    // =========================================================================
    task automatic run_simple_loop_test();
        $display("\n=============================================================");
        $display("Simple Loop Test - Verify branch behavior");
        $display("=============================================================\n");
        
        // Load simple loop program
        instruction_mem[0] = 32'h00000293;  // addi    t0, x0, 0
        instruction_mem[1] = 32'h00A00313;  // addi    t1, x0, 10
        instruction_mem[2] = 32'h00000393;  // addi    t2, x0, 0
        instruction_mem[3] = 32'h00138393;  // addi    t2, t2, 1
        instruction_mem[4] = 32'h00128293;  // addi    t0, t0, 1
        instruction_mem[5] = 32'hFE62CCE3;  // blt     t0, t1, -8
        instruction_mem[6] = 32'h00502023;  // sw      t0, 0(x0)
        instruction_mem[7] = 32'h00602223;  // sw      t1, 4(x0)
        instruction_mem[8] = 32'h00702423;  // sw      t2, 8(x0)
        instruction_mem[9] = 32'h00000013;  // nop
        
        // Clear data memory
        for (int i = 0; i < 16; i++) data_mem[i] = 0;
        
        rst = 1'b1;
        #20;
        rst = 1'b0;
        
        // Wait for loop to complete (10 iterations * ~5 cycles each + overhead)
        #1000;
        
        // Verify results
        $display("Results:");
        $display("  t0 (counter) = %0d (expected 10)", data_mem[0]);
        $display("  t1 (limit)   = %0d (expected 10)", data_mem[1]);
        $display("  t2 (accum)   = %0d (expected 10)", data_mem[2]);
        
        if (data_mem[0] == 10 && data_mem[1] == 10 && data_mem[2] == 10) begin
            $display("PASS: Simple loop test passed!");
            checked += 3;
        end else begin
            $display("FAIL: Simple loop test failed!");
            checked += 3;
            errors += 3;
        end
    endtask

    // =========================================================================
    // Main Test Sequence
    // =========================================================================
    initial begin
        // VCD dump for waveform analysis
        $dumpfile("tb_chacha20.vcd");
        $dumpvars(0, tb_chacha20);
        
        // Initialize
        checked = 0;
        errors = 0;
        
        $display("=============================================================");
        $display("    ChaCha20 Full Block Testbench");
        $display("=============================================================\n");
        
        // First, run simple loop test to verify branch works
        run_simple_loop_test();
        
        // Load test vector and program
        load_chacha20_test_vector();
        load_chacha20_program();
        
        $display("\nInput state (ChaCha20 constants + key + counter + nonce):");
        for (int i = 0; i < 16; i++) begin
            $display("  state[%2d] = 0x%08X", i, data_mem[i]);
        end
        
        // Reset and run
        rst = 1'b1;
        #20;
        rst = 1'b0;
        
        $display("\nRunning ChaCha20 block (20 rounds = 10 double-rounds)...");
        $display("This executes ~3500 instructions with heavy ROL usage.\n");
        
        // Wait for completion (10 rounds @ ~1.3ms each = ~13ms, add margin)
        #20000000;
        
        // =====================
        // Verify Results
        // =====================
        $display("=============================================================");
        $display("Verifying ChaCha20 results...");
        $display("=============================================================\n");
        
        // Check round counter (should be 10, stored at 0x200 = word 128)
        if (data_mem[128] == 32'd10) begin
            $display("PASS: Completed 10 double-rounds (counter = %d)", data_mem[128]);
            checked++;
        end else begin
            $display("FAIL: Round counter expected 10, got %d", data_mem[128]);
            checked++;
            errors++;
        end
        
        // Check CPOP integrity (stored at 0x204 = word 129)
        if (data_mem[129] > 0 && data_mem[129] <= 32) begin
            $display("PASS: CPOP integrity check = %d bits", data_mem[129]);
            checked++;
        end else begin
            $display("FAIL: CPOP expected 1-32, got %d", data_mem[129]);
            checked++;
            errors++;
        end
        
        // Check that output differs from input (output at 0x40 = word 16)
        $display("\nOutput state (after 20 rounds):");
        for (int i = 0; i < 16; i++) begin
            $display("  output[%2d] = 0x%08X", i, data_mem[16 + i]);
            
            // Verify output changed from input
            if (data_mem[16 + i] != data_mem[i]) begin
                checked++;
            end else begin
                $display("    WARNING: output[%d] unchanged from input!", i);
                checked++;
                errors++;
            end
        end
        
        // =====================
        // Summary
        // =====================
        $display("\n=============================================================");
        $display("                      Test Summary");
        $display("=============================================================");
        $display("  Total Checks: %0d", checked);
        $display("  Passed:       %0d", checked - errors);
        $display("  Failed:       %0d", errors);
        $display("=============================================================\n");
        
        if (errors) begin
            display_fail();
        end else begin
            display_pass();
        end
        
        $finish;
    end

endmodule

